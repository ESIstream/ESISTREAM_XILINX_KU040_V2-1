-------------------------------------------------------------------------------
-- This is free and unencumbered software released into the public domain.
--
-- Anyone is free to copy, modify, publish, use, compile, sell, or distribute
-- this software, either in source code form or as a compiled bitstream, for 
-- any purpose, commercial or non-commercial, and by any means.
--
-- In jurisdictions that recognize copyright laws, the author or authors of 
-- this software dedicate any and all copyright interest in the software to 
-- the public domain. We make this dedication for the benefit of the public at
-- large and to the detriment of our heirs and successors. We intend this 
-- dedication to be an overt act of relinquishment in perpetuity of all present
-- and future rights to this software under copyright law.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR 
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN 
-- ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION
-- WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
--
-- THIS DISCLAIMER MUST BE RETAINED AS PART OF THIS FILE AT ALL TIMES. 
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity edge_detect is
  generic (
    EDGE_TYPE : string := "RISING"
    );
  port (
    clk           : in  std_logic;
    din           : in  std_logic;
    edge_detected : out std_logic
    );
end edge_detect;

architecture rtl of edge_detect is

  signal din_t : std_logic := '0';
  signal din_r : std_logic_vector(1 downto 0) := (others => '0');

begin

  din_t <= din;

  din_reg : process (clk)
  begin
    if rising_edge (clk) then
      din_r(0) <= din_t;
      din_r(1) <= din_r(0);
    end if;
  end process;

  rising_edge_detect : if EDGE_TYPE = "RISING" generate
  begin
    process (clk)
    begin
      if rising_edge (clk) then
        edge_detected <= din_r(0) and (not din_r(1));
      end if;
    end process;
  end generate;

  falling_edge_detect : if EDGE_TYPE = "FALLING" generate
  begin
    process (clk)
    begin
      if rising_edge (clk) then
        edge_detected <= din_r(1) and (not din_r(0));
      end if;
    end process;
  end generate;

end architecture rtl;
